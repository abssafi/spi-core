package wb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    `include "wb_packet.sv"

endpackage