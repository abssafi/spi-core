class wb_master_monitor extends superClass;
    function new();
        
    endfunction //new()
endclass //wb_master_monitor extends superClass